module  sva_imm_test;

endmodule
